
module boot_code
(
    input  logic        CLK,
    input  logic        RSTN,

    input  logic        CSN,
    input  logic [9:0]  A,
    output logic [31:0] Q
  );

  const logic [0:899] [31:0] mem = {
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h0100006F,
    32'h0100006F,
    32'h0080006F,
    32'h0040006F,
    32'h0000006F,
    32'h00000093,
    32'h81868106,
    32'h82868206,
    32'h83868306,
    32'h84868406,
    32'h85868506,
    32'h86868606,
    32'h87868706,
    32'h88868806,
    32'h89868906,
    32'h8A868A06,
    32'h8B868B06,
    32'h8C868C06,
    32'h8D868D06,
    32'h8E868E06,
    32'h8F868F06,
    32'h20000117,
    32'hF3010113,
    32'h00000D17,
    32'h618D0D13,
    32'h00000D97,
    32'h610D8D93,
    32'h01BD5763,
    32'h000D2023,
    32'hDDE30D11,
    32'h0513FFAD,
    32'h05930000,
    32'h00EF0000,
    32'h00000140,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h11010000,
<<<<<<< HEAD
    32'h03100593,
    32'hCE064501,
    32'hCA26CC22,
    32'hC64EC84A,
    32'hC256C452,
    32'h1F6000EF,
    32'h50000737,
    32'hAAAA16B7,
    32'h869387BA,
    32'hA22B1116,
    32'h26B700D7,
    32'h8693BBBB,
    32'hC3942226,
    32'hCCCC36B7,
    32'h33368693,
    32'h46B7C714,
    32'h8693DDDD,
    32'hC7544446,
    32'hEEEE56B7,
    32'h002DC7B7,
    32'h55568693,
    32'h6C078793,
    32'hC0FBCB14,
    32'h00010037,
    32'h09B70001,
    32'h49255000,
    32'h002DCAB7,
    32'h01498A13,
    32'h0049A48B,
    32'hD7B34471,
    32'hB7B34084,
    32'h1471F647,
    32'h05778513,
    32'h00F96463,
    32'h03078513,
    32'h20C000EF,
    32'hFFC433E3,
    32'h00EF4529,
    32'h87932020,
    32'hC0FB6C0A,
    32'h00010037,
    32'h95E30001,
    32'h0537FD49,
    32'h45D10001,
    32'h3D450513,
    32'h19E000EF,
    32'h00010537,
    32'h03900593,
    32'h3EC50513,
    32'h18E000EF,
    32'h00010537,
    32'h03800593,
    32'h42850513,
    32'h17E000EF,
    32'h00010537,
    32'h03800593,
    32'h46450513,
    32'h16E000EF,
    32'h00010537,
    32'h03800593,
    32'h4A050513,
    32'h15E000EF,
    32'h00010537,
    32'h03800593,
    32'h4DC50513,
    32'h14E000EF,
    32'h00010537,
    32'h03800593,
    32'h51850513,
    32'h13E000EF,
    32'h00010537,
    32'h03800593,
    32'h55450513,
    32'h12E000EF,
    32'h00010537,
    32'h03700593,
    32'h59050513,
    32'h11E000EF,
    32'h00010537,
    32'h03800593,
    32'h5C850513,
    32'h10E000EF,
    32'h166000EF,
    32'h87936785,
    32'hC0FBBB87,
    32'h00010037,
    32'h05370001,
    32'h05930001,
    32'h05130230,
    32'h00EF6045,
    32'h00EF0EC0,
    32'h45291440,
    32'h128000EF,
=======
    32'h450145E1,
    32'hCC22CE06,
    32'hC84ACA26,
    32'hC452C64E,
    32'h00EFC256,
    32'h00EF1FA0,
    32'h07372AA0,
    32'h16B72200,
    32'h87BAAAAA,
    32'h11168693,
    32'h00D7A22B,
    32'hBBBB26B7,
    32'h22268693,
    32'h36B7C394,
    32'h8693CCCC,
    32'hC7143336,
    32'hDDDD46B7,
    32'h44468693,
    32'h56B7C754,
    32'hC7B7EEEE,
    32'h8693002D,
    32'h87935556,
    32'hCB146C07,
    32'h0037C0FB,
    32'h00010001,
    32'h220009B7,
    32'hCAB74925,
    32'h8A13002D,
    32'hA48B0149,
    32'h44710049,
    32'h4084D7B3,
    32'hF647B7B3,
    32'h85131471,
    32'h64630577,
    32'h851300F9,
    32'h00EF0307,
    32'h33E320C0,
    32'h4529FFC4,
    32'h202000EF,
    32'h6C0A8793,
    32'h0037C0FB,
    32'h00010001,
    32'hFD4995E3,
    32'h00010537,
    32'h051345D1,
    32'h00EF4485,
    32'h053719E0,
    32'h05930001,
    32'h05130390,
    32'h00EF4605,
    32'h053718E0,
    32'h05930001,
    32'h05130380,
    32'h00EF49C5,
    32'h053717E0,
    32'h05930001,
    32'h05130380,
    32'h00EF4D85,
    32'h053716E0,
    32'h05930001,
    32'h05130380,
    32'h00EF5145,
    32'h053715E0,
    32'h05930001,
    32'h05130380,
    32'h00EF5505,
    32'h053714E0,
    32'h05930001,
    32'h05130380,
    32'h00EF58C5,
    32'h053713E0,
    32'h05930001,
    32'h05130380,
    32'h00EF5C85,
    32'h053712E0,
    32'h05930001,
    32'h05130370,
    32'h00EF6045,
    32'h053711E0,
    32'h05930001,
    32'h05130380,
    32'h00EF63C5,
    32'h00EF10E0,
    32'h67851660,
    32'hBB878793,
    32'h0037C0FB,
    32'h00010001,
    32'h00010537,
    32'h02300593,
    32'h67850513,
    32'h0EC000EF,
    32'h144000EF,
    32'h00EF4529,
    32'h44611280,
    32'h00EF4481,
    32'h15331060,
    32'h14610085,
    32'h3AE38CC9,
    32'hAB63FF84,
    32'h446103F4,
    32'h00EF4901,
    32'h15330EE0,
    32'h14610085,
    32'h00A96933,
    32'hFF8439E3,
    32'h0124A023,
>>>>>>> b6f7552f80b2d3c0291eeeb705874daf8e7b2fe6
    32'h44814461,
    32'h0D4000EF,
    32'h00851533,
    32'h8CC91461,
    32'hFF843AE3,
<<<<<<< HEAD
    32'h03F4AB63,
    32'h49014461,
    32'h0EE000EF,
    32'h00851533,
    32'h69331461,
    32'h39E300A9,
    32'hA023FF84,
    32'h44610124,
    32'h00EF4481,
    32'h15330D40,
    32'h14610085,
    32'h3AE38CC9,
    32'hB9E3FF84,
    32'h0537FDF4,
    32'h05130001,
    32'h45956285,
    32'h08A000EF,
    32'h00010537,
    32'h051345ED,
    32'h00EF6305,
    32'h00EF07C0,
    32'h07B70D40,
    32'h67375000,
    32'hC71C1A10,
    32'h08078793,
    32'h00078067,
=======
    32'hFDF4B9E3,
    32'h00010537,
    32'h69C50513,
    32'h00EF4595,
    32'h053708A0,
    32'h45ED0001,
    32'h6A450513,
    32'h07C000EF,
    32'h0D4000EF,
    32'h260007B7,
    32'h1A106737,
    32'h8793C71C,
    32'h80670807,
    32'h00010007,
>>>>>>> b6f7552f80b2d3c0291eeeb705874daf8e7b2fe6
    32'h00010001,
    32'h450140F2,
    32'h44D24462,
    32'h49B24942,
    32'h4A924A22,
    32'h80826105,
    32'h1A106737,
    32'h43100711,
    32'h1A1007B7,
    32'hC0164633,
    32'h8693C310,
    32'h85130047,
    32'hD81300C7,
    32'h07130085,
    32'hF5930830,
    32'hC1180FF5,
    32'h0106A023,
    32'h0A700713,
    32'h00B7A42B,
    32'h478DC398,
    32'h429CC11C,
    32'h0F07F793,
    32'hC017C7B3,
    32'h8082C29C,
    32'h1A100737,
    32'hC1850751,
    32'h04000693,
    32'hF793431C,
    32'hDFED0207,
    32'h0015460B,
    32'h1A1007B7,
    32'hC39015FD,
    32'hE29916FD,
    32'h8082F1F5,
    32'h8082F1F5,
    32'h1A100737,
    32'h431C0751,
    32'hFC17B7B3,
    32'h07B7DFED,
    32'h43881A10,
    32'h0FF57513,
    32'h07378082,
    32'h07511A10,
    32'hF793431C,
<<<<<<< HEAD
    32'hDFED0407,
=======
    32'hDFED0207,
    32'h1A1007B7,
    32'h8082C388,
    32'h1A100737,
    32'h431C0751,
    32'h0407F793,
    32'h8082DFED,
    32'h280006B7,
    32'h429C06C1,
    32'h28000737,
    32'h00779613,
    32'hFE065BE3,
    32'h0ADFA7B7,
    32'h00470613,
    32'h6A678793,
    32'h17B7C21C,
    32'h06930017,
    32'h87930087,
    32'h0731E207,
    32'h431CC29C,
    32'hC007C7B3,
    32'h6785C31C,
    32'hBB878793,
    32'h0037C0FB,
    32'h00010001,
    32'h8793678D,
    32'h07373A87,
    32'hC31C2800,
    32'h12C1D0FB,
    32'h00010001,
    32'h879367C1,
    32'h07374107,
    32'hCB1C2800,
    32'h0641D0FB,
    32'h00010001,
>>>>>>> b6f7552f80b2d3c0291eeeb705874daf8e7b2fe6
    32'h00008082,
    32'h20202020,
    32'h20202020,
    32'h20202020,
    32'h20202020,
    32'h0A555520,
    32'h00000000,
    32'h20202020,
    32'h20202020,
    32'h20202020,
    32'h55555555,
    32'h55555555,
    32'h55555555,
    32'h20202020,
    32'h55552020,
    32'h55555555,
    32'h55555555,
    32'h20202020,
    32'h55555555,
    32'h55202055,
    32'h55555555,
    32'h0000000A,
    32'h20202020,
    32'h20202020,
    32'h55202020,
    32'h20205555,
    32'h20555520,
    32'h55552020,
    32'h20202055,
    32'h20202020,
    32'h20202055,
    32'h55202020,
    32'h20202055,
    32'h20205520,
    32'h20202020,
    32'h0A552020,
    32'h00000000,
    32'h20202020,
    32'h20202020,
    32'h55552020,
    32'h20202055,
    32'h20555520,
    32'h55202020,
    32'h20205555,
    32'h20202020,
    32'h20202055,
    32'h55202020,
    32'h20202020,
    32'h20205520,
    32'h20202020,
    32'h0A552020,
    32'h00000000,
    32'h20202020,
    32'h20202020,
    32'h55552020,
    32'h20202020,
    32'h20555520,
    32'h20202020,
    32'h20205555,
    32'h20202020,
    32'h55555555,
    32'h20205555,
    32'h20202020,
    32'h20205520,
    32'h20202020,
    32'h0A552020,
    32'h00000000,
    32'h20202020,
    32'h20202020,
    32'h55552020,
    32'h20202020,
    32'h20555520,
    32'h55202020,
    32'h20205555,
    32'h20202020,
    32'h20202055,
    32'h20202020,
    32'h20544F49,
    32'h20205520,
    32'h20202020,
    32'h0A552020,
    32'h00000000,
    32'h20202020,
    32'h20202020,
    32'h55202020,
    32'h55555555,
    32'h20555520,
    32'h55555555,
    32'h20202020,
    32'h20202020,
    32'h20202055,
    32'h49412020,
    32'h20202020,
    32'h20205520,
    32'h20202020,
    32'h0A552020,
    32'h00000000,
    32'h20202020,
    32'h20202020,
    32'h20202020,
    32'h55552020,
    32'h55555555,
    32'h20205555,
    32'h20202020,
    32'h20202020,
    32'h20202055,
    32'h20202020,
    32'h20202020,
    32'h20555520,
    32'h20202020,
    32'h0A555520,
    32'h00000000,
    32'h20202020,
    32'h20202020,
    32'h20202020,
    32'h20202020,
    32'h20555555,
    32'h52202020,
    32'h2D435349,
    32'h20202056,
    32'h20202055,
    32'h43202020,
    32'h20706968,
    32'h55552020,
    32'h20202020,
    32'h000A5555,
    32'h20202020,
    32'h20202020,
    32'h20202020,
    32'h55202020,
    32'h55555555,
    32'h20202020,
    32'h20202020,
    32'h55552020,
    32'h55555555,
    32'h20202055,
    32'h20202020,
    32'h55202020,
    32'h55555555,
    32'h0A0A0A55,
    32'h00000000,
    32'h61656C50,
    32'h55206573,
    32'h616F6C70,
    32'h72502064,
    32'h6172676F,
    32'h6976206D,
    32'h41552061,
    32'h2E205452,
    32'h000A2E2E,
    32'h656E6F44,
    32'h0000000A,
    32'h706D754A,
    32'h20676E69,
    32'h49206F74,
    32'h7274736E,
    32'h69746375,
    32'h52206E6F,
    32'h000A4D41,
    32'h00000010,
    32'h00000000,
    32'h00527A01,
    32'h01010401,
    32'h00020D1B,
    32'h00000028,
    32'h00000018,
<<<<<<< HEAD
    32'hFFFFFAAA,
    32'h0000020C,
=======
    32'hFFFFFA36,
    32'h0000020E,
>>>>>>> b6f7552f80b2d3c0291eeeb705874daf8e7b2fe6
    32'h200E4200,
    32'h7F011152,
    32'h117E0811,
    32'h12117D09,
    32'h7B13117C,
    32'h117A1411,
    32'h00007915,
    32'h00000010,
    32'h00000044,
<<<<<<< HEAD
    32'hFFFFFC8A,
=======
    32'hFFFFFC18,
>>>>>>> b6f7552f80b2d3c0291eeeb705874daf8e7b2fe6
    32'h00000048,
    32'h00000000,
    32'h00000010,
    32'h00000058,
<<<<<<< HEAD
    32'hFFFFFCBE,
=======
    32'hFFFFFC4C,
>>>>>>> b6f7552f80b2d3c0291eeeb705874daf8e7b2fe6
    32'h0000002C,
    32'h00000000,
    32'h00000010,
    32'h0000006C,
<<<<<<< HEAD
    32'hFFFFFCD6,
=======
    32'hFFFFFC64,
>>>>>>> b6f7552f80b2d3c0291eeeb705874daf8e7b2fe6
    32'h0000001A,
    32'h00000000,
    32'h00000010,
    32'h00000080,
<<<<<<< HEAD
    32'hFFFFFCDC,
=======
    32'hFFFFFC6A,
>>>>>>> b6f7552f80b2d3c0291eeeb705874daf8e7b2fe6
    32'h00000016,
    32'h00000000,
    32'h00000010,
    32'h00000094,
<<<<<<< HEAD
    32'hFFFFFCDE,
    32'h00000010,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
=======
    32'hFFFFFC6C,
    32'h00000010,
    32'h00000000,
    32'h00000010,
    32'h000000A8,
    32'hFFFFFC68,
    32'h00000072,
>>>>>>> b6f7552f80b2d3c0291eeeb705874daf8e7b2fe6
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000};

  logic [9:0] A_Q;

  always_ff @(posedge CLK, negedge RSTN)
  begin
    if (~RSTN)
      A_Q <= '0;
    else
      if (~CSN)
        A_Q <= A;
  end

  assign Q = mem[A_Q];

endmodule