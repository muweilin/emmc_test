
module boot_code0
(
    input  logic        CLK,
    input  logic        RSTN,

    input  logic        CSN,
    input  logic [9:0]  A,
    output logic [31:0] Q
  );

  const logic [0:547] [31:0] mem = {
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h0100006F,
    32'h0100006F,
    32'h0080006F,
    32'h0040006F,
    32'h0000006F,
    32'h00000093,
    32'h81868106,
    32'h82868206,
    32'h83868306,
    32'h84868406,
    32'h85868506,
    32'h86868606,
    32'h87868706,
    32'h88868806,
    32'h89868906,
    32'h8A868A06,
    32'h8B868B06,
    32'h8C868C06,
    32'h8D868D06,
    32'h8E868E06,
    32'h8F868F06,
    32'h00100117,
    32'hF3010113,
    32'h00000D17,
    32'h670D0D13,
    32'h00000D97,
    32'h668D8D93,
    32'h01BD5763,
    32'h000D2023,
    32'hDDE30D11,
    32'h0513FFAD,
    32'h05930000,
    32'h00EF0000,
    32'h00000140,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h11410000,
    32'h03100593,
    32'hC6064501,
    32'hC226C422,
    32'h00EFC04A,
    32'h85371A20,
    32'h45D90000,
    32'h36450513,
    32'h1DC000EF,
    32'h00008537,
    32'h051345D1,
    32'h00EF37C5,
    32'h85371CE0,
    32'h45D10000,
    32'h39450513,
    32'h1C0000EF,
    32'h00008537,
    32'h03900593,
    32'h3AC50513,
    32'h1B0000EF,
    32'h00008537,
    32'h03800593,
    32'h3E850513,
    32'h1A0000EF,
    32'h00008537,
    32'h03800593,
    32'h42450513,
    32'h190000EF,
    32'h00008537,
    32'h03800593,
    32'h46050513,
    32'h180000EF,
    32'h00008537,
    32'h03800593,
    32'h49C50513,
    32'h170000EF,
    32'h00008537,
    32'h03800593,
    32'h4D850513,
    32'h160000EF,
    32'h00008537,
    32'h03800593,
    32'h51450513,
    32'h150000EF,
    32'h00008537,
    32'h03800593,
    32'h55050513,
    32'h140000EF,
    32'h00008537,
    32'h03800593,
    32'h58C50513,
    32'h130000EF,
    32'h00008537,
    32'h03800593,
    32'h5C850513,
    32'h120000EF,
    32'h00008537,
    32'h03700593,
    32'h60450513,
    32'h110000EF,
    32'h00008537,
    32'h03800593,
    32'h63C50513,
    32'h100000EF,
    32'h142000EF,
    32'h87936785,
    32'hC0FBBB87,
    32'h00010037,
    32'h85370001,
    32'h05930000,
    32'h05130230,
    32'h00EF6785,
    32'h44610DE0,
    32'h11E000EF,
    32'h00EF4481,
    32'h15330FE0,
    32'h14610085,
    32'h3AE38CC9,
    32'hAB63FF84,
    32'h446103F4,
    32'h00EF4901,
    32'h15330E60,
    32'h14610085,
    32'h00A96933,
    32'hFF8439E3,
    32'h0124A023,
    32'h44814461,
    32'h0CC000EF,
    32'h00851533,
    32'h8CC91461,
    32'hFF843AE3,
    32'hFDF4B9E3,
    32'h00008537,
    32'h69C50513,
    32'h00EF4595,
    32'h85370820,
    32'h45ED0000,
    32'h6A450513,
    32'h074000EF,
    32'h0B6000EF,
    32'h1A1067B7,
    32'h0007A423,
    32'h08000793,
    32'h00078067,
    32'h00010001,
    32'h40B20001,
    32'h44224501,
    32'h49024492,
    32'h80820141,
    32'h1A106737,
    32'h43100711,
    32'h1A1007B7,
    32'hC0164633,
    32'h8693C310,
    32'h85130047,
    32'hD81300C7,
    32'h07130085,
    32'hF5930830,
    32'hC1180FF5,
    32'h0106A023,
    32'h0A700713,
    32'h00B7A42B,
    32'h478DC398,
    32'h429CC11C,
    32'h0F07F793,
    32'hC017C7B3,
    32'h8082C29C,
    32'h1A100737,
    32'hC1850751,
    32'h04000693,
    32'hF793431C,
    32'hDFED0207,
    32'h0015460B,
    32'h1A1007B7,
    32'hC39015FD,
    32'hE29916FD,
    32'h8082F1F5,
    32'h8082F1F5,
    32'h1A100737,
    32'h431C0751,
    32'hFC17B7B3,
    32'h07B7DFED,
    32'h43881A10,
    32'h0FF57513,
    32'h07378082,
    32'h07511A10,
    32'hF793431C,
    32'hDFED0407,
    32'h00008082,
    32'h20202020,
    32'h20202020,
    32'h20202020,
    32'h55552020,
    32'h55555555,
    32'h00000A55,
    32'h20202020,
    32'h20202020,
    32'h20202020,
    32'h20202020,
    32'h0A555555,
    32'h00000000,
    32'h20202020,
    32'h20202020,
    32'h20202020,
    32'h20202020,
    32'h0A555520,
    32'h00000000,
    32'h20202020,
    32'h20202020,
    32'h20202020,
    32'h55555555,
    32'h55555555,
    32'h55555555,
    32'h20202020,
    32'h55552020,
    32'h55555555,
    32'h55555555,
    32'h20202020,
    32'h55555555,
    32'h55202055,
    32'h55555555,
    32'h0000000A,
    32'h20202020,
    32'h20202020,
    32'h55202020,
    32'h20205555,
    32'h20555520,
    32'h55552020,
    32'h20202055,
    32'h20202020,
    32'h20202055,
    32'h55202020,
    32'h20202055,
    32'h20205520,
    32'h20202020,
    32'h0A552020,
    32'h00000000,
    32'h20202020,
    32'h20202020,
    32'h55552020,
    32'h20202055,
    32'h20555520,
    32'h55202020,
    32'h20205555,
    32'h20202020,
    32'h20202055,
    32'h20202020,
    32'h20202055,
    32'h20205520,
    32'h20202020,
    32'h0A552020,
    32'h00000000,
    32'h20202020,
    32'h20202020,
    32'h55555520,
    32'h20202020,
    32'h20555520,
    32'h20202020,
    32'h20555555,
    32'h20202020,
    32'h20202055,
    32'h55202020,
    32'h20202020,
    32'h20205520,
    32'h20202020,
    32'h0A552020,
    32'h00000000,
    32'h20202020,
    32'h20202020,
    32'h55555520,
    32'h20202020,
    32'h20555520,
    32'h20202020,
    32'h20555555,
    32'h20202020,
    32'h20202055,
    32'h20552020,
    32'h20202020,
    32'h20205520,
    32'h20202020,
    32'h0A552020,
    32'h00000000,
    32'h20202020,
    32'h20202020,
    32'h55555520,
    32'h20202020,
    32'h20555520,
    32'h20202020,
    32'h20555555,
    32'h20202020,
    32'h55555555,
    32'h20205555,
    32'h20202020,
    32'h20205520,
    32'h20202020,
    32'h0A552020,
    32'h00000000,
    32'h20202020,
    32'h20202020,
    32'h55552020,
    32'h20202020,
    32'h20555520,
    32'h55202020,
    32'h20205555,
    32'h20202020,
    32'h20202055,
    32'h20202020,
    32'h20544F49,
    32'h20205520,
    32'h20202020,
    32'h0A552020,
    32'h00000000,
    32'h20202020,
    32'h20202020,
    32'h55552020,
    32'h20202055,
    32'h20555520,
    32'h55552020,
    32'h20202055,
    32'h20202020,
    32'h20202055,
    32'h20202020,
    32'h20202020,
    32'h20205520,
    32'h20202020,
    32'h0A552020,
    32'h00000000,
    32'h20202020,
    32'h20202020,
    32'h55202020,
    32'h55555555,
    32'h20555520,
    32'h55555555,
    32'h20202020,
    32'h20202020,
    32'h20202055,
    32'h49412020,
    32'h20202020,
    32'h20205520,
    32'h20202020,
    32'h0A552020,
    32'h00000000,
    32'h20202020,
    32'h20202020,
    32'h20202020,
    32'h55552020,
    32'h55555555,
    32'h20205555,
    32'h20202020,
    32'h20202020,
    32'h20202055,
    32'h20202020,
    32'h20202020,
    32'h20555520,
    32'h20202020,
    32'h0A555520,
    32'h00000000,
    32'h20202020,
    32'h20202020,
    32'h20202020,
    32'h20202020,
    32'h20555555,
    32'h52202020,
    32'h2D435349,
    32'h20202056,
    32'h20202055,
    32'h43202020,
    32'h20706968,
    32'h55552020,
    32'h20202020,
    32'h000A5555,
    32'h20202020,
    32'h20202020,
    32'h20202020,
    32'h55202020,
    32'h55555555,
    32'h20202020,
    32'h20202020,
    32'h55552020,
    32'h55555555,
    32'h20202055,
    32'h20202020,
    32'h55202020,
    32'h55555555,
    32'h0A0A0A55,
    32'h00000000,
    32'h61656C50,
    32'h55206573,
    32'h616F6C70,
    32'h72502064,
    32'h6172676F,
    32'h6976206D,
    32'h41552061,
    32'h2E205452,
    32'h000A2E2E,
    32'h656E6F44,
    32'h0000000A,
    32'h706D754A,
    32'h20676E69,
    32'h49206F74,
    32'h7274736E,
    32'h69746375,
    32'h52206E6F,
    32'h000A4D41,
    32'h00000010,
    32'h00000000,
    32'h00527A01,
    32'h01010401,
    32'h00020D1B,
    32'h00000020,
    32'h00000018,
    32'hFFFFFA36,
    32'h000001B2,
    32'h100E4200,
    32'h7F01114E,
    32'h117E0811,
    32'h12117D09,
    32'h0000007C,
    32'h00000010,
    32'h0000003C,
    32'hFFFFFBC4,
    32'h00000048,
    32'h00000000,
    32'h00000010,
    32'h00000050,
    32'hFFFFFBF8,
    32'h0000002C,
    32'h00000000,
    32'h00000010,
    32'h00000064,
    32'hFFFFFC10,
    32'h0000001A,
    32'h00000000,
    32'h00000010,
    32'h00000078,
    32'hFFFFFC16,
    32'h00000010,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000};

  logic [9:0] A_Q;

  always_ff @(posedge CLK, negedge RSTN)
  begin
    if (~RSTN)
      A_Q <= '0;
    else
      if (~CSN)
        A_Q <= A;
  end

  assign Q = mem[A_Q];

endmodule