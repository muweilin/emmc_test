
module boot_code
(
    input  logic        CLK,
    input  logic        RSTN,

    input  logic        CSN,
    input  logic [9:0]  A,
    output logic [31:0] Q
  );

  const logic [0:899] [31:0] mem = {
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h0100006F,
    32'h0100006F,
    32'h0080006F,
    32'h0040006F,
    32'h0000006F,
    32'h00000093,
    32'h81868106,
    32'h82868206,
    32'h83868306,
    32'h84868406,
    32'h85868506,
    32'h86868606,
    32'h87868706,
    32'h88868806,
    32'h89868906,
    32'h8A868A06,
    32'h8B868B06,
    32'h8C868C06,
    32'h8D868D06,
    32'h8E868E06,
    32'h8F868F06,
    32'h52FF4117,
    32'hF3010113,
    32'h00000D17,
    32'h618D0D13,
    32'h00000D97,
    32'h610D8D93,
    32'h01BD5763,
    32'h000D2023,
    32'hDDE30D11,
    32'h0513FFAD,
    32'h05930000,
    32'h00EF0000,
    32'h00000140,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h11010000,
    32'h03100593,
    32'hCE064501,
    32'hCA26CC22,
    32'hC64EC84A,
    32'hC256C452,
    32'h1F6000EF,
    32'h50000737,
    32'hAAAA16B7,
    32'h869387BA,
    32'hA22B1116,
    32'h26B700D7,
    32'h8693BBBB,
    32'hC3942226,
    32'hCCCC36B7,
    32'h33368693,
    32'h46B7C714,
    32'h8693DDDD,
    32'hC7544446,
    32'hEEEE56B7,
    32'h002DC7B7,
    32'h55568693,
    32'h6C078793,
    32'hC0FBCB14,
    32'h00010037,
    32'h09B70001,
    32'h49255000,
    32'h002DCAB7,
    32'h01498A13,
    32'h0049A48B,
    32'hD7B34471,
    32'hB7B34084,
    32'h1471F647,
    32'h05778513,
    32'h00F96463,
    32'h03078513,
    32'h20C000EF,
    32'hFFC433E3,
    32'h00EF4529,
    32'h87932020,
    32'hC0FB6C0A,
    32'h00010037,
    32'h95E30001,
    32'h0537FD49,
    32'h45D10001,
    32'h3D450513,
    32'h19E000EF,
    32'h00010537,
    32'h03900593,
    32'h3EC50513,
    32'h18E000EF,
    32'h00010537,
    32'h03800593,
    32'h42850513,
    32'h17E000EF,
    32'h00010537,
    32'h03800593,
    32'h46450513,
    32'h16E000EF,
    32'h00010537,
    32'h03800593,
    32'h4A050513,
    32'h15E000EF,
    32'h00010537,
    32'h03800593,
    32'h4DC50513,
    32'h14E000EF,
    32'h00010537,
    32'h03800593,
    32'h51850513,
    32'h13E000EF,
    32'h00010537,
    32'h03800593,
    32'h55450513,
    32'h12E000EF,
    32'h00010537,
    32'h03700593,
    32'h59050513,
    32'h11E000EF,
    32'h00010537,
    32'h03800593,
    32'h5C850513,
    32'h10E000EF,
    32'h166000EF,
    32'h87936785,
    32'hC0FBBB87,
    32'h00010037,
    32'h05370001,
    32'h05930001,
    32'h05130230,
    32'h00EF6045,
    32'h00EF0EC0,
    32'h45291440,
    32'h128000EF,
    32'h44814461,
    32'h106000EF,
    32'h00851533,
    32'h8CC91461,
    32'hFF843AE3,
    32'h03F4AB63,
    32'h49014461,
    32'h0EE000EF,
    32'h00851533,
    32'h69331461,
    32'h39E300A9,
    32'hA023FF84,
    32'h44610124,
    32'h00EF4481,
    32'h15330D40,
    32'h14610085,
    32'h3AE38CC9,
    32'hB9E3FF84,
    32'h0537FDF4,
    32'h05130001,
    32'h45956285,
    32'h08A000EF,
    32'h00010537,
    32'h051345ED,
    32'h00EF6305,
    32'h00EF07C0,
    32'h07B70D40,
    32'h67375000,
    32'hC71C1A10,
    32'h08078793,
    32'h00078067,
    32'h00010001,
    32'h40F20001,
    32'h44624501,
    32'h494244D2,
    32'h4A2249B2,
    32'h61054A92,
    32'h67378082,
    32'h07111A10,
    32'h07B74310,
    32'h46331A10,
    32'hC310C016,
    32'h00478693,
    32'h00C78513,
    32'h0085D813,
    32'h08300713,
    32'h0FF5F593,
    32'hA023C118,
    32'h07130106,
    32'hA42B0A70,
    32'hC39800B7,
    32'hC11C478D,
    32'hF793429C,
    32'hC7B30F07,
    32'hC29CC017,
    32'h07378082,
    32'h07511A10,
    32'h0693C185,
    32'h431C0400,
    32'h0207F793,
    32'h460BDFED,
    32'h07B70015,
    32'h15FD1A10,
    32'h16FDC390,
    32'hF1F5E299,
    32'hF1F58082,
    32'h07378082,
    32'h07511A10,
    32'hB7B3431C,
    32'hDFEDFC17,
    32'h1A1007B7,
    32'h75134388,
    32'h80820FF5,
    32'h1A100737,
    32'h431C0751,
    32'h0207F793,
    32'h07B7DFED,
    32'hC3881A10,
    32'h07378082,
    32'h07511A10,
    32'hF793431C,
    32'hDFED0407,
    32'h00008082,
    32'h20202020,
    32'h20202020,
    32'h20202020,
    32'h20202020,
    32'h0A555520,
    32'h00000000,
    32'h20202020,
    32'h20202020,
    32'h20202020,
    32'h55555555,
    32'h55555555,
    32'h55555555,
    32'h20202020,
    32'h55552020,
    32'h55555555,
    32'h55555555,
    32'h20202020,
    32'h55555555,
    32'h55202055,
    32'h55555555,
    32'h0000000A,
    32'h20202020,
    32'h20202020,
    32'h55202020,
    32'h20205555,
    32'h20555520,
    32'h55552020,
    32'h20202055,
    32'h20202020,
    32'h20202055,
    32'h55202020,
    32'h20202055,
    32'h20205520,
    32'h20202020,
    32'h0A552020,
    32'h00000000,
    32'h20202020,
    32'h20202020,
    32'h55552020,
    32'h20202055,
    32'h20555520,
    32'h55202020,
    32'h20205555,
    32'h20202020,
    32'h20202055,
    32'h55202020,
    32'h20202020,
    32'h20205520,
    32'h20202020,
    32'h0A552020,
    32'h00000000,
    32'h20202020,
    32'h20202020,
    32'h55552020,
    32'h20202020,
    32'h20555520,
    32'h20202020,
    32'h20205555,
    32'h20202020,
    32'h55555555,
    32'h20205555,
    32'h20202020,
    32'h20205520,
    32'h20202020,
    32'h0A552020,
    32'h00000000,
    32'h20202020,
    32'h20202020,
    32'h55552020,
    32'h20202020,
    32'h20555520,
    32'h55202020,
    32'h20205555,
    32'h20202020,
    32'h20202055,
    32'h20202020,
    32'h20544F49,
    32'h20205520,
    32'h20202020,
    32'h0A552020,
    32'h00000000,
    32'h20202020,
    32'h20202020,
    32'h55202020,
    32'h55555555,
    32'h20555520,
    32'h55555555,
    32'h20202020,
    32'h20202020,
    32'h20202055,
    32'h49412020,
    32'h20202020,
    32'h20205520,
    32'h20202020,
    32'h0A552020,
    32'h00000000,
    32'h20202020,
    32'h20202020,
    32'h20202020,
    32'h55552020,
    32'h55555555,
    32'h20205555,
    32'h20202020,
    32'h20202020,
    32'h20202055,
    32'h20202020,
    32'h20202020,
    32'h20555520,
    32'h20202020,
    32'h0A555520,
    32'h00000000,
    32'h20202020,
    32'h20202020,
    32'h20202020,
    32'h20202020,
    32'h20555555,
    32'h52202020,
    32'h2D435349,
    32'h20202056,
    32'h20202055,
    32'h43202020,
    32'h20706968,
    32'h55552020,
    32'h20202020,
    32'h000A5555,
    32'h20202020,
    32'h20202020,
    32'h20202020,
    32'h55202020,
    32'h55555555,
    32'h20202020,
    32'h20202020,
    32'h55552020,
    32'h55555555,
    32'h20202055,
    32'h20202020,
    32'h55202020,
    32'h55555555,
    32'h0A0A0A55,
    32'h00000000,
    32'h61656C50,
    32'h55206573,
    32'h616F6C70,
    32'h72502064,
    32'h6172676F,
    32'h6976206D,
    32'h41552061,
    32'h2E205452,
    32'h000A2E2E,
    32'h656E6F44,
    32'h0000000A,
    32'h706D754A,
    32'h20676E69,
    32'h49206F74,
    32'h7274736E,
    32'h69746375,
    32'h52206E6F,
    32'h000A4D41,
    32'h00000010,
    32'h00000000,
    32'h00527A01,
    32'h01010401,
    32'h00020D1B,
    32'h00000028,
    32'h00000018,
    32'hFFFFFAAA,
    32'h0000020C,
    32'h200E4200,
    32'h7F011154,
    32'h117E0811,
    32'h12117D09,
    32'h7B13117C,
    32'h117A1411,
    32'h00007915,
    32'h00000010,
    32'h00000044,
    32'hFFFFFC8A,
    32'h00000048,
    32'h00000000,
    32'h00000010,
    32'h00000058,
    32'hFFFFFCBE,
    32'h0000002C,
    32'h00000000,
    32'h00000010,
    32'h0000006C,
    32'hFFFFFCD6,
    32'h0000001A,
    32'h00000000,
    32'h00000010,
    32'h00000080,
    32'hFFFFFCDC,
    32'h00000016,
    32'h00000000,
    32'h00000010,
    32'h00000094,
    32'hFFFFFCDE,
    32'h00000010,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000};

  logic [9:0] A_Q;

  always_ff @(posedge CLK, negedge RSTN)
  begin
    if (~RSTN)
      A_Q <= '0;
    else
      if (~CSN)
        A_Q <= A;
  end

  assign Q = mem[A_Q];

endmodule