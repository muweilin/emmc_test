
module boot_code
(
    input  logic        CLK,
    input  logic        RSTN,

    input  logic        CSN,
    input  logic [9:0]  A,
    output logic [31:0] Q
  );

  const logic [0:899] [31:0] mem = {
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h0100006F,
    32'h0100006F,
    32'h0080006F,
    32'h0040006F,
    32'h0000006F,
    32'h00000093,
    32'h81868106,
    32'h82868206,
    32'h83868306,
    32'h84868406,
    32'h85868506,
    32'h86868606,
    32'h87868706,
    32'h88868806,
    32'h89868906,
    32'h8A868A06,
    32'h8B868B06,
    32'h8C868C06,
    32'h8D868D06,
    32'h8E868E06,
    32'h8F868F06,
    32'h52FF4117,
    32'hF3010113,
    32'h00001D17,
    32'h8D8D0D13,
    32'h00001D97,
    32'h8D0D8D93,
    32'h01BD5763,
    32'h000D2023,
    32'hDDE30D11,
    32'h0513FFAD,
    32'h05930000,
    32'h00EF0000,
    32'h00000140,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h715D0000,
    32'h03100593,
    32'hC6864501,
    32'hC2A6C4A2,
    32'hDE4EC0CA,
    32'hDA56DC52,
    32'hD65ED85A,
    32'hD266D462,
    32'h00EFD06A,
    32'h47113EC0,
    32'h1A1027B7,
    32'h00010537,
    32'h45F5C3D8,
    32'h5A450513,
    32'h41E000EF,
    32'h00010537,
    32'h051345D1,
    32'h00EF5C45,
    32'h05374100,
    32'h05930001,
    32'h05130390,
    32'h00EF5DC5,
    32'h05374000,
    32'h05930001,
    32'h05130380,
    32'h00EF6185,
    32'h05373F00,
    32'h05930001,
    32'h05130380,
    32'h00EF6545,
    32'h05373E00,
    32'h05930001,
    32'h05130380,
    32'h00EF6905,
    32'h05373D00,
    32'h05930001,
    32'h05130380,
    32'h00EF6CC5,
    32'h05373C00,
    32'h05930001,
    32'h05130380,
    32'h00EF7085,
    32'h05373B00,
    32'h05930001,
    32'h05130380,
    32'h00EF7445,
    32'h05373A00,
    32'h05930001,
    32'h05130370,
    32'h00EF7805,
    32'h05373900,
    32'h05930001,
    32'h05130380,
    32'h00EF7B85,
    32'h00EF3800,
    32'h46813A80,
    32'h45A14601,
    32'h09F00513,
    32'h240000EF,
    32'h45014581,
    32'h26C000EF,
    32'h02000513,
    32'h274000EF,
    32'h45014581,
    32'h28C000EF,
    32'h02000593,
    32'h00EF0028,
    32'h27B72B40,
    32'h47220120,
    32'h84D78793,
    32'h02F70163,
    32'h010227B7,
    32'h94D78793,
    32'h00F70B63,
    32'h00010537,
    32'h02400593,
    32'h7F450513,
    32'h322000EF,
    32'h0693A001,
    32'h46010200,
    32'h454D45A1,
    32'h1E4000EF,
    32'h0A000513,
    32'h220000EF,
    32'h45014581,
    32'h238000EF,
    32'h0A000593,
    32'h00EF0068,
    32'h4BC22600,
    32'h44524962,
    32'h8B5E4A32,
    32'h4AF289CA,
    32'h1BF42363,
    32'h00011537,
    32'h051345F5,
    32'h00EF8485,
    32'h00EF2D80,
    32'h15373000,
    32'h45C50001,
    32'h86850513,
    32'h2C6000EF,
    32'h2EE000EF,
    32'h41F45793,
    32'h0167D493,
    32'h00940733,
    32'hEAA7B7B3,
    32'hEAA73733,
    32'h1487A45B,
    32'h409704B3,
    32'h04805363,
    32'h4C018B52,
    32'h414B8D33,
    32'h865A6C85,
    32'h02000693,
    32'h454D45A1,
    32'h15C000EF,
    32'h00EF6521,
    32'h458119A0,
    32'h00EF4501,
    32'h0C051B20,
    32'h016D0533,
    32'h00EF65A1,
    32'h9B661D80,
    32'hFD841BE3,
    32'h00C41793,
    32'h00FB8B33,
    32'h06939A3E,
    32'h86520200,
    32'h454D45A1,
    32'h00549413,
    32'h120000EF,
    32'h00EF8522,
    32'h458115E0,
    32'h00EF4501,
    32'h85A21760,
    32'h00EF855A,
    32'h00EF1A00,
    32'h553318C0,
    32'h3CE31005,
    32'h1537FE15,
    32'h45C50001,
    32'h87C50513,
    32'h21E000EF,
    32'h246000EF,
    32'h41FAD793,
    32'h0167D693,
    32'h00DA8733,
    32'hEAA7B7B3,
    32'h3733048A,
    32'hA45BEAA7,
    32'h94D21557,
    32'h40D70A33,
    32'h04805263,
    32'h4A8189A6,
    32'h40990BB3,
    32'h864E6B05,
    32'h02000693,
    32'h454D45A1,
    32'h0B0000EF,
    32'h00EF6521,
    32'h45810EE0,
    32'h00EF4501,
    32'h0A851060,
    32'h013B8533,
    32'h00EF65A1,
    32'h99DA12C0,
    32'hFD541BE3,
    32'h09B30432,
    32'h94A20089,
    32'h02000693,
    32'h45A18626,
    32'h005A1413,
    32'h00EF454D,
    32'h85220760,
    32'h0B4000EF,
    32'h45014581,
    32'h0CC000EF,
    32'h854E85A2,
    32'h0F6000EF,
    32'h00011537,
    32'h051345E9,
    32'h00EF8905,
    32'h00EF1800,
    32'h67B71A80,
    32'hA4231A10,
    32'h07B70007,
    32'h87935000,
    32'h80670807,
    32'h00010007,
    32'h00010001,
    32'h450140B6,
    32'h44964426,
    32'h59F24906,
    32'h5AD25A62,
    32'h5BB25B42,
    32'h5C925C22,
    32'h61615D02,
    32'h15378082,
    32'h05930001,
    32'h05130290,
    32'h00EF81C5,
    32'hA0011340,
    32'h08136811,
    32'h06A2F008,
    32'h02000713,
    32'h1A1027B7,
    32'hF6B38F0D,
    32'hB5B30106,
    32'h1533F265,
    32'h881300E5,
    32'h87130087,
    32'h8DD500C7,
    32'h202307C1,
    32'hC31000A8,
    32'h8082C38C,
    32'h553305C2,
    32'h8DC91005,
    32'h1A1027B7,
    32'h8082CBCC,
    32'h1A102737,
    32'h431C0741,
    32'hC63E1141,
    32'hD7B347B2,
    32'h05421007,
    32'hC62A8D5D,
    32'hC31C47B2,
    32'h80820141,
    32'h05A14785,
    32'h00B795B3,
    32'h00A79533,
    32'h87936785,
    32'h8DFDF007,
    32'hEE853533,
    32'h27B78D4D,
    32'hC3881A10,
    32'h27B78082,
    32'h439C1A10,
    32'hC63E1141,
    32'h01414532,
    32'h97B38082,
    32'h1141D455,
    32'hF455B5B3,
    32'hC581C43E,
    32'h078547A2,
    32'hC602C43E,
    32'h273746B2,
    32'h47A21A10,
    32'h02070813,
    32'h02F6D563,
    32'h97B3431C,
    32'hDFEDCF07,
    32'h258347B2,
    32'h46B20008,
    32'hC6360685,
    32'h078A0810,
    32'hFFC62603,
    32'h67A346A2,
    32'h4FE300B5,
    32'h0141FCD6,
    32'h67378082,
    32'h07111A10,
    32'h07B74310,
    32'h46331A10,
    32'hC310C016,
    32'h00478693,
    32'h00C78513,
    32'h0085D813,
    32'h08300713,
    32'h0FF5F593,
    32'hA023C118,
    32'h07130106,
    32'hA42B0A70,
    32'hC39800B7,
    32'hC11C478D,
    32'hF793429C,
    32'hC7B30F07,
    32'hC29CC017,
    32'h07378082,
    32'h07511A10,
    32'h0693C185,
    32'h431C0400,
    32'h0207F793,
    32'h460BDFED,
    32'h07B70015,
    32'h15FD1A10,
    32'h16FDC390,
    32'hF1F5E299,
    32'hF1F58082,
    32'h07378082,
    32'h07511A10,
    32'hF793431C,
    32'hDFED0407,
    32'h00008082,
    32'h72617453,
    32'h676E6974,
    32'h50755720,
    32'h302E3175,
    32'h524F4320,
    32'h2E2E2045,
    32'h2E2E2E2E,
    32'h0000000A,
    32'h20202020,
    32'h20202020,
    32'h20202020,
    32'h20202020,
    32'h0A555520,
    32'h00000000,
    32'h20202020,
    32'h20202020,
    32'h20202020,
    32'h55555555,
    32'h55555555,
    32'h55555555,
    32'h20202020,
    32'h55552020,
    32'h55555555,
    32'h55555555,
    32'h20202020,
    32'h55555555,
    32'h55202055,
    32'h55555555,
    32'h0000000A,
    32'h20202020,
    32'h20202020,
    32'h55202020,
    32'h20205555,
    32'h20555520,
    32'h55552020,
    32'h20202055,
    32'h20202020,
    32'h20202055,
    32'h55202020,
    32'h20202055,
    32'h20205520,
    32'h20202020,
    32'h0A552020,
    32'h00000000,
    32'h20202020,
    32'h20202020,
    32'h55552020,
    32'h20202055,
    32'h20555520,
    32'h55202020,
    32'h20205555,
    32'h20202020,
    32'h20202055,
    32'h55202020,
    32'h20202020,
    32'h20205520,
    32'h20202020,
    32'h0A552020,
    32'h00000000,
    32'h20202020,
    32'h20202020,
    32'h55552020,
    32'h20202020,
    32'h20555520,
    32'h20202020,
    32'h20205555,
    32'h20202020,
    32'h55555555,
    32'h20205555,
    32'h20202020,
    32'h20205520,
    32'h20202020,
    32'h0A552020,
    32'h00000000,
    32'h20202020,
    32'h20202020,
    32'h55552020,
    32'h20202020,
    32'h20555520,
    32'h55202020,
    32'h20205555,
    32'h20202020,
    32'h20202055,
    32'h20202020,
    32'h20544F49,
    32'h20205520,
    32'h20202020,
    32'h0A552020,
    32'h00000000,
    32'h20202020,
    32'h20202020,
    32'h55202020,
    32'h55555555,
    32'h20555520,
    32'h55555555,
    32'h20202020,
    32'h20202020,
    32'h20202055,
    32'h49412020,
    32'h20202020,
    32'h20205520,
    32'h20202020,
    32'h0A552020,
    32'h00000000,
    32'h20202020,
    32'h20202020,
    32'h20202020,
    32'h55552020,
    32'h55555555,
    32'h20205555,
    32'h20202020,
    32'h20202020,
    32'h20202055,
    32'h20202020,
    32'h20202020,
    32'h20555520,
    32'h20202020,
    32'h0A555520,
    32'h00000000,
    32'h20202020,
    32'h20202020,
    32'h20202020,
    32'h20202020,
    32'h20555555,
    32'h52202020,
    32'h2D435349,
    32'h20202056,
    32'h20202055,
    32'h43202020,
    32'h20706968,
    32'h55552020,
    32'h20202020,
    32'h000A5555,
    32'h20202020,
    32'h20202020,
    32'h20202020,
    32'h55202020,
    32'h55555555,
    32'h20202020,
    32'h20202020,
    32'h55552020,
    32'h55555555,
    32'h20202055,
    32'h20202020,
    32'h55202020,
    32'h55555555,
    32'h0A0A0A55,
    32'h00000000,
    32'h4F525245,
    32'h53203A52,
    32'h736E6170,
    32'h206E6F69,
    32'h20495053,
    32'h73616C66,
    32'h6F6E2068,
    32'h6F662074,
    32'h0A646E75,
    32'h00000000,
    32'h4F525245,
    32'h54203A52,
    32'h65726568,
    32'h20736920,
    32'h70206F6E,
    32'h72676F72,
    32'h69206D61,
    32'h6F79206E,
    32'h66207275,
    32'h6873616C,
    32'h0000000A,
    32'h64616F4C,
    32'h20676E69,
    32'h67616D69,
    32'h72662065,
    32'h53206D6F,
    32'h66204950,
    32'h6873616C,
    32'h0000000A,
    32'h64616F4C,
    32'h20676E69,
    32'h65646F63,
    32'h2E2E2E20,
    32'h0000000A,
    32'h64616F4C,
    32'h20676E69,
    32'h61746164,
    32'h2E2E2E20,
    32'h0000000A,
    32'h706D754A,
    32'h20676E69,
    32'h75206F74,
    32'h20726573,
    32'h67616D69,
    32'h2E2E2065,
    32'h00000A2E,
    32'h00000010,
    32'h00000000,
    32'h00527A01,
    32'h01010401,
    32'h00020D1B,
    32'h00000038,
    32'h00000018,
    32'hFFFFF84A,
    32'h00000326,
    32'h500E4200,
    32'h7F01115E,
    32'h117E0811,
    32'h12117D09,
    32'h7B13117C,
    32'h117A1411,
    32'h16117915,
    32'h77171178,
    32'h11761811,
    32'h1A117519,
    32'h00000074,
    32'h00000010,
    32'h00000054,
    32'hFFFFFB34,
    32'h00000034,
    32'h00000000,
    32'h00000010,
    32'h00000068,
    32'hFFFFFB54,
    32'h00000010,
    32'h00000000,
    32'h00000010,
    32'h0000007C,
    32'hFFFFFB50,
    32'h00000020,
    32'h100E4A00,
    32'h00000010,
    32'h00000090,
    32'hFFFFFB5C,
    32'h00000022,
    32'h00000000,
    32'h00000010,
    32'h000000A4,
    32'hFFFFFB6A,
    32'h00000010,
    32'h100E4800,
    32'h00000010,
    32'h000000B8,
    32'hFFFFFB66,
    32'h00000050,
    32'h100E4600,
    32'h00000010,
    32'h000000CC,
    32'hFFFFFBA2,
    32'h00000048,
    32'h00000000,
    32'h00000010,
    32'h000000E0,
    32'hFFFFFBD6,
    32'h0000002C,
    32'h00000000,
    32'h00000010,
    32'h000000F4,
    32'hFFFFFBEE,
    32'h00000010,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000};

  logic [9:0] A_Q;

  always_ff @(posedge CLK, negedge RSTN)
  begin
    if (~RSTN)
      A_Q <= '0;
    else
      if (~CSN)
        A_Q <= A;
  end

  assign Q = mem[A_Q];

endmodule